`timescale 1ns/1ps

module FIR_TwoParallel (
    input  logic clk,
    input  logic rst,
    input  logic signed [15:0] in_even,
    input  logic signed [15:0] in_odd,
    output logic signed [63:0] out_even,
    output logic signed [63:0] out_odd
);

    parameter int NUM_TAPS = 102;
    localparam int HALF_TAPS = NUM_TAPS / 2;

    // Coefficient memory (fixed)
    localparam logic signed [31:0] coeffs [NUM_TAPS-1:0] = '{
        32'b11111111111110000101000100011100,
        32'b11111111111000110010100001001110,
        32'b11111111101101000000010001110011,
        32'b11111111010111011101110000111000,
        32'b11111110110101011110110010000100,
        32'b11111110000110010100100000001110,
        32'b11111101001100100110001111000010,
        32'b11111100001111001011001111010110,
        32'b11111011011001000010101110010000,
        32'b11111010110111110010101000110100,
        32'b11111010111000101110000110111000,
        32'b11111011100101000100011110011001,
        32'b11111100111110010111010100010101,
        32'b11111110111100000101010000001000,
        32'b00000001001011101110100110110101,
        32'b00000011010011110110001000001100,
        32'b00000100111001101000100110000110,
        32'b00000101100111111010111100110001,
        32'b00000101010101100010100111100101,
        32'b00000100001001000010111110000001,
        32'b00000010011000001101001000111111,
        32'b00000000100010111001101111101100,
        32'b11111111001010100000100110100001,
        32'b11111110101000000110001000011001,
        32'b11111111000100011111011111101110,
        32'b00000000010100111100110110111100,
        32'b00000001111101110111111000010001,
        32'b00000011011011001011111111100001,
        32'b00000100001100000000101100011010,
        32'b00000011111101111001110010001101,
        32'b00000010110011110110100011111110,
        32'b00000001000110010010100000101101,
        32'b11111111011011100111010000000100,
        32'b11111110011011010011001101101110,
        32'b11111110011111101100110010101111,
        32'b11111111101011011100101000111111,
        32'b00000001100110100010000111100001,
        32'b00000011100100101110100110111001,
        32'b00000100110011111011100110100011,
        32'b00000100101110000110100000111010,
        32'b00000011001000110110001101011100,
        32'b00000000011101000010001100100101,
        32'b11111101100011000100010101000111,
        32'b11111011100100000011000000011100,
        32'b11111011100011110001010101110010,
        32'b11111110001010001101000101110100,
        32'b00000011010011101001110010101011,
        32'b00001010001101001001100110000011,
        32'b00010001011110111100101000011100,
        32'b00010111100010100111010001011110,
        32'b00011010111110100000001110101110,
        32'b00011010111110100000001110101110,
        32'b00010111100010100111010001011110,
        32'b00010001011110111100101000011100,
        32'b00001010001101001001100110000011,
        32'b00000011010011101001110010101011,
        32'b11111110001010001101000101110100,
        32'b11111011100011110001010101110010,
        32'b11111011100100000011000000011100,
        32'b11111101100011000100010101000111,
        32'b00000000011101000010001100100101,
        32'b00000011001000110110001101011100,
        32'b00000100101110000110100000111010,
        32'b00000100110011111011100110100011,
        32'b00000011100100101110100110111001,
        32'b00000001100110100010000111100001,
        32'b11111111101011011100101000111111,
        32'b11111110011111101100110010101111,
        32'b11111110011011010011001101101110,
        32'b11111111011011100111010000000100,
        32'b00000001000110010010100000101101,
        32'b00000010110011110110100011111110,
        32'b00000011111101111001110010001101,
        32'b00000100001100000000101100011010,
        32'b00000011011011001011111111100001,
        32'b00000001111101110111111000010001,
        32'b00000000010100111100110110111100,
        32'b11111111000100011111011111101110,
        32'b11111110101000000110001000011001,
        32'b11111111001010100000100110100001,
        32'b00000000100010111001101111101100,
        32'b00000010011000001101001000111111,
        32'b00000100001001000010111110000001,
        32'b00000101010101100010100111100101,
        32'b00000101100111111010111100110001,
        32'b00000100111001101000100110000110,
        32'b00000011010011110110001000001100,
        32'b00000001001011101110100110110101,
        32'b11111110111100000101010000001000,
        32'b11111100111110010111010100010101,
        32'b11111011100101000100011110011001,
        32'b11111010111000101110000110111000,
        32'b11111010110111110010101000110100,
        32'b11111011011001000010101110010000,
        32'b11111100001111001011001111010110,
        32'b11111101001100100110001111000010,
        32'b11111110000110010100100000001110,
        32'b11111110110101011110110010000100,
        32'b11111111010111011101110000111000,
        32'b11111111101101000000010001110011,
        32'b11111111111000110010100001001110,
        32'b11111111111110000101000100011100
    };
  // Internal delay lines for even/odd indexed inputs
    logic signed [15:0] delay_even [HALF_TAPS-1:0];
    logic signed [15:0] delay_odd  [HALF_TAPS-1:0];

    // Intermediate sums
    logic signed [63:0] accum_even, accum_odd, accum_combined;
    logic signed [63:0] prev_odd_sum;

    // Shift registers and state
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            prev_odd_sum <= 0;
            for (int k = 0; k < HALF_TAPS; k++) begin
                delay_even[k] <= 0;
                delay_odd[k]  <= 0;
            end
        end else begin
            for (int k = HALF_TAPS-1; k > 0; k--) begin
                delay_even[k] <= delay_even[k-1];
                delay_odd[k]  <= delay_odd[k-1];
            end
            delay_even[0] <= in_even;
            delay_odd[0]  <= in_odd;
            prev_odd_sum <= accum_odd;
        end
    end

    // FIR multiply-accumulate logic
    always_comb begin
        accum_even     = 0;
        accum_odd      = 0;
        accum_combined = 0;

        for (int k = 0; k < HALF_TAPS; k++) begin
            accum_even     += delay_even[k] * coeffs[2*k];
            accum_odd      += delay_odd[k]  * coeffs[2*k+1];
            accum_combined += (delay_even[k] + delay_odd[k]) * 
                              (coeffs[2*k] + coeffs[2*k+1]);
        end
    end

    // Final output assignment with scaling
    assign out_even = (accum_even + prev_odd_sum) >>> 31;
    assign out_odd  = (accum_combined - accum_even - accum_odd) >>> 31;

endmodule
