`timescale 1ns/1ps

module three_parallel_pipeline (
    input  logic              clk,         // Master clock
    input  logic              rst,         // Asynchronous reset
    input  logic signed [15:0] d_in,       // Single input sample
    output logic signed [63:0] d_out       // Filtered output
);

    // Overall number of FIR taps
    parameter int NUM_TAPS = 102;

    // Stored coefficients (scaled Q1.31 format)
        localparam logic signed [31:0] coef [TAPS-1:0] = '{
        32'b11111111111110000101000100011100,
        32'b11111111111000110010100001001110,
        32'b11111111101101000000010001110011,
        32'b11111111010111011101110000111000,
        32'b11111110110101011110110010000100,
        32'b11111110000110010100100000001110,
        32'b11111101001100100110001111000010,
        32'b11111100001111001011001111010110,
        32'b11111011011001000010101110010000,
        32'b11111010110111110010101000110100,
        32'b11111010111000101110000110111000,
        32'b11111011100101000100011110011001,
        32'b11111100111110010111010100010101,
        32'b11111110111100000101010000001000,
        32'b00000001001011101110100110110101,
        32'b00000011010011110110001000001100,
        32'b00000100111001101000100110000110,
        32'b00000101100111111010111100110001,
        32'b00000101010101100010100111100101,
        32'b00000100001001000010111110000001,
        32'b00000010011000001101001000111111,
        32'b00000000100010111001101111101100,
        32'b11111111001010100000100110100001,
        32'b11111110101000000110001000011001,
        32'b11111111000100011111011111101110,
        32'b00000000010100111100110110111100,
        32'b00000001111101110111111000010001,
        32'b00000011011011001011111111100001,
        32'b00000100001100000000101100011010,
        32'b00000011111101111001110010001101,
        32'b00000010110011110110100011111110,
        32'b00000001000110010010100000101101,
        32'b11111111011011100111010000000100,
        32'b11111110011011010011001101101110,
        32'b11111110011111101100110010101111,
        32'b11111111101011011100101000111111,
        32'b00000001100110100010000111100001,
        32'b00000011100100101110100110111001,
        32'b00000100110011111011100110100011,
        32'b00000100101110000110100000111010,
        32'b00000011001000110110001101011100,
        32'b00000000011101000010001100100101,
        32'b11111101100011000100010101000111,
        32'b11111011100100000011000000011100,
        32'b11111011100011110001010101110010,
        32'b11111110001010001101000101110100,
        32'b00000011010011101001110010101011,
        32'b00001010001101001001100110000011,
        32'b00010001011110111100101000011100,
        32'b00010111100010100111010001011110,
        32'b00011010111110100000001110101110,
        32'b00011010111110100000001110101110,
        32'b00010111100010100111010001011110,
        32'b00010001011110111100101000011100,
        32'b00001010001101001001100110000011,
        32'b00000011010011101001110010101011,
        32'b11111110001010001101000101110100,
        32'b11111011100011110001010101110010,
        32'b11111011100100000011000000011100,
        32'b11111101100011000100010101000111,
        32'b00000000011101000010001100100101,
        32'b00000011001000110110001101011100,
        32'b00000100101110000110100000111010,
        32'b00000100110011111011100110100011,
        32'b00000011100100101110100110111001,
        32'b00000001100110100010000111100001,
        32'b11111111101011011100101000111111,
        32'b11111110011111101100110010101111,
        32'b11111110011011010011001101101110,
        32'b11111111011011100111010000000100,
        32'b00000001000110010010100000101101,
        32'b00000010110011110110100011111110,
        32'b00000011111101111001110010001101,
        32'b00000100001100000000101100011010,
        32'b00000011011011001011111111100001,
        32'b00000001111101110111111000010001,
        32'b00000000010100111100110110111100,
        32'b11111111000100011111011111101110,
        32'b11111110101000000110001000011001,
        32'b11111111001010100000100110100001,
        32'b00000000100010111001101111101100,
        32'b00000010011000001101001000111111,
        32'b00000100001001000010111110000001,
        32'b00000101010101100010100111100101,
        32'b00000101100111111010111100110001,
        32'b00000100111001101000100110000110,
        32'b00000011010011110110001000001100,
        32'b00000001001011101110100110110101,
        32'b11111110111100000101010000001000,
        32'b11111100111110010111010100010101,
        32'b11111011100101000100011110011001,
        32'b11111010111000101110000110111000,
        32'b11111010110111110010101000110100,
        32'b11111011011001000010101110010000,
        32'b11111100001111001011001111010110,
        32'b11111101001100100110001111000010,
        32'b11111110000110010100100000001110,
        32'b11111110110101011110110010000100,
        32'b11111111010111011101110000111000,
        32'b11111111101101000000010001110011,
        32'b11111111111000110010100001001110,
        32'b11111111111110000101000100011100
    };
     // Delay line sized for pipeline logic
    // (One sample per clock but extended storage for partial accumulation)
    logic signed [15:0] shift_buffer [2*NUM_TAPS-2:0];
    
    // Pipeline for accumulate
    logic signed [63:0] accum_stage [NUM_TAPS-1:0];

    // Shift samples on each rising edge or reset
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            for (int i = 0; i < 2*NUM_TAPS-1; i++) begin
                shift_buffer[i] <= 16'sd0;
            end
        end else begin
            for (int i = 2*NUM_TAPS-2; i > 0; i--) begin
                shift_buffer[i] <= shift_buffer[i - 1];
            end
            // Insert the latest input sample
            shift_buffer[0] <= d_in;
        end
    end

    // Accumulate partial products in pipeline stages
    always_ff @(posedge clk) begin
        accum_stage[0] <= d_in * coeff_mem[0];
        for (int k = 1; k < NUM_TAPS; k++) begin
            accum_stage[k] <= accum_stage[k-1] 
                              + shift_buffer[2*(k-1)+1] * coeff_mem[k];
        end
    end

    // Shift right by 31 bits to align final Q1.31 product
    assign d_out = accum_stage[NUM_TAPS-1] >>> 31;

endmodule
